`define Psum_BITS 24 


